module clock_buf (out,in);

output out;
input in;

buf G1(out,in);

endmodule